`ifndef definitions_SVH
`define definitions_SVH
                                
`define OPCODE_I_TYPE      7'b00?0011
`define OPCODE_I_JALR_TYPE 7'b1100111
`define OPCODE_S_TYPE      7'b0100011
`define OPCODE_B_TYPE      7'b1100011
`define OPCODE_U_TYPE      7'b0?10111
`define OPCODE_J_TYPE      7'b1101111

`endif // definitions_SVH
