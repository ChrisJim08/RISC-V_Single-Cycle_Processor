'timescale 1ns / 1ps

module flopr();


endmodule