'timescale 1ns / 1ps

module alu();


endmodule