'timescale 1ns / 1ps

module alu_controller ();


endmodule